library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity power_lut_8 is
port(
    clk_i:in std_logic;
    a: in std_logic_vector(7 downto 0);
    z: out unsigned(15 downto 0)
);
end power_lut_8;
architecture rtl of power_lut_8 is
begin
    power_lut:process(clk_i)
    begin
        if rising_edge(clk_i) then
            case a is
                when "00000000" => z <= "0000000000000000";
                when "00000001" => z <= "0000000000000001";
                when "00000010" => z <= "0000000000000100";
                when "00000011" => z <= "0000000000001001";
                when "00000100" => z <= "0000000000010000";
                when "00000101" => z <= "0000000000011001";
                when "00000110" => z <= "0000000000100100";
                when "00000111" => z <= "0000000000110001";
                when "00001000" => z <= "0000000001000000";
                when "00001001" => z <= "0000000001010001";
                when "00001010" => z <= "0000000001100100";
                when "00001011" => z <= "0000000001111001";
                when "00001100" => z <= "0000000010010000";
                when "00001101" => z <= "0000000010101001";
                when "00001110" => z <= "0000000011000100";
                when "00001111" => z <= "0000000011100001";
                when "00010000" => z <= "0000000100000000";
                when "00010001" => z <= "0000000100100001";
                when "00010010" => z <= "0000000101000100";
                when "00010011" => z <= "0000000101101001";
                when "00010100" => z <= "0000000110010000";
                when "00010101" => z <= "0000000110111001";
                when "00010110" => z <= "0000000111100100";
                when "00010111" => z <= "0000001000010001";
                when "00011000" => z <= "0000001001000000";
                when "00011001" => z <= "0000001001110001";
                when "00011010" => z <= "0000001010100100";
                when "00011011" => z <= "0000001011011001";
                when "00011100" => z <= "0000001100010000";
                when "00011101" => z <= "0000001101001001";
                when "00011110" => z <= "0000001110000100";
                when "00011111" => z <= "0000001111000001";
                when "00100000" => z <= "0000010000000000";
                when "00100001" => z <= "0000010001000001";
                when "00100010" => z <= "0000010010000100";
                when "00100011" => z <= "0000010011001001";
                when "00100100" => z <= "0000010100010000";
                when "00100101" => z <= "0000010101011001";
                when "00100110" => z <= "0000010110100100";
                when "00100111" => z <= "0000010111110001";
                when "00101000" => z <= "0000011001000000";
                when "00101001" => z <= "0000011010010001";
                when "00101010" => z <= "0000011011100100";
                when "00101011" => z <= "0000011100111001";
                when "00101100" => z <= "0000011110010000";
                when "00101101" => z <= "0000011111101001";
                when "00101110" => z <= "0000100001000100";
                when "00101111" => z <= "0000100010100001";
                when "00110000" => z <= "0000100100000000";
                when "00110001" => z <= "0000100101100001";
                when "00110010" => z <= "0000100111000100";
                when "00110011" => z <= "0000101000101001";
                when "00110100" => z <= "0000101010010000";
                when "00110101" => z <= "0000101011111001";
                when "00110110" => z <= "0000101101100100";
                when "00110111" => z <= "0000101111010001";
                when "00111000" => z <= "0000110001000000";
                when "00111001" => z <= "0000110010110001";
                when "00111010" => z <= "0000110100100100";
                when "00111011" => z <= "0000110110011001";
                when "00111100" => z <= "0000111000010000";
                when "00111101" => z <= "0000111010001001";
                when "00111110" => z <= "0000111100000100";
                when "00111111" => z <= "0000111110000001";
                when "01000000" => z <= "0001000000000000";
                when "01000001" => z <= "0001000010000001";
                when "01000010" => z <= "0001000100000100";
                when "01000011" => z <= "0001000110001001";
                when "01000100" => z <= "0001001000010000";
                when "01000101" => z <= "0001001010011001";
                when "01000110" => z <= "0001001100100100";
                when "01000111" => z <= "0001001110110001";
                when "01001000" => z <= "0001010001000000";
                when "01001001" => z <= "0001010011010001";
                when "01001010" => z <= "0001010101100100";
                when "01001011" => z <= "0001010111111001";
                when "01001100" => z <= "0001011010010000";
                when "01001101" => z <= "0001011100101001";
                when "01001110" => z <= "0001011111000100";
                when "01001111" => z <= "0001100001100001";
                when "01010000" => z <= "0001100100000000";
                when "01010001" => z <= "0001100110100001";
                when "01010010" => z <= "0001101001000100";
                when "01010011" => z <= "0001101011101001";
                when "01010100" => z <= "0001101110010000";
                when "01010101" => z <= "0001110000111001";
                when "01010110" => z <= "0001110011100100";
                when "01010111" => z <= "0001110110010001";
                when "01011000" => z <= "0001111001000000";
                when "01011001" => z <= "0001111011110001";
                when "01011010" => z <= "0001111110100100";
                when "01011011" => z <= "0010000001011001";
                when "01011100" => z <= "0010000100010000";
                when "01011101" => z <= "0010000111001001";
                when "01011110" => z <= "0010001010000100";
                when "01011111" => z <= "0010001101000001";
                when "01100000" => z <= "0010010000000000";
                when "01100001" => z <= "0010010011000001";
                when "01100010" => z <= "0010010110000100";
                when "01100011" => z <= "0010011001001001";
                when "01100100" => z <= "0010011100010000";
                when "01100101" => z <= "0010011111011001";
                when "01100110" => z <= "0010100010100100";
                when "01100111" => z <= "0010100101110001";
                when "01101000" => z <= "0010101001000000";
                when "01101001" => z <= "0010101100010001";
                when "01101010" => z <= "0010101111100100";
                when "01101011" => z <= "0010110010111001";
                when "01101100" => z <= "0010110110010000";
                when "01101101" => z <= "0010111001101001";
                when "01101110" => z <= "0010111101000100";
                when "01101111" => z <= "0011000000100001";
                when "01110000" => z <= "0011000100000000";
                when "01110001" => z <= "0011000111100001";
                when "01110010" => z <= "0011001011000100";
                when "01110011" => z <= "0011001110101001";
                when "01110100" => z <= "0011010010010000";
                when "01110101" => z <= "0011010101111001";
                when "01110110" => z <= "0011011001100100";
                when "01110111" => z <= "0011011101010001";
                when "01111000" => z <= "0011100001000000";
                when "01111001" => z <= "0011100100110001";
                when "01111010" => z <= "0011101000100100";
                when "01111011" => z <= "0011101100011001";
                when "01111100" => z <= "0011110000010000";
                when "01111101" => z <= "0011110100001001";
                when "01111110" => z <= "0011111000000100";
                when "01111111" => z <= "0011111100000001";
                when "10000000" => z <= "0100000000000000";
                when "10000001" => z <= "0011111100000001";
                when "10000010" => z <= "0011111000000100";
                when "10000011" => z <= "0011110100001001";
                when "10000100" => z <= "0011110000010000";
                when "10000101" => z <= "0011101100011001";
                when "10000110" => z <= "0011101000100100";
                when "10000111" => z <= "0011100100110001";
                when "10001000" => z <= "0011100001000000";
                when "10001001" => z <= "0011011101010001";
                when "10001010" => z <= "0011011001100100";
                when "10001011" => z <= "0011010101111001";
                when "10001100" => z <= "0011010010010000";
                when "10001101" => z <= "0011001110101001";
                when "10001110" => z <= "0011001011000100";
                when "10001111" => z <= "0011000111100001";
                when "10010000" => z <= "0011000100000000";
                when "10010001" => z <= "0011000000100001";
                when "10010010" => z <= "0010111101000100";
                when "10010011" => z <= "0010111001101001";
                when "10010100" => z <= "0010110110010000";
                when "10010101" => z <= "0010110010111001";
                when "10010110" => z <= "0010101111100100";
                when "10010111" => z <= "0010101100010001";
                when "10011000" => z <= "0010101001000000";
                when "10011001" => z <= "0010100101110001";
                when "10011010" => z <= "0010100010100100";
                when "10011011" => z <= "0010011111011001";
                when "10011100" => z <= "0010011100010000";
                when "10011101" => z <= "0010011001001001";
                when "10011110" => z <= "0010010110000100";
                when "10011111" => z <= "0010010011000001";
                when "10100000" => z <= "0010010000000000";
                when "10100001" => z <= "0010001101000001";
                when "10100010" => z <= "0010001010000100";
                when "10100011" => z <= "0010000111001001";
                when "10100100" => z <= "0010000100010000";
                when "10100101" => z <= "0010000001011001";
                when "10100110" => z <= "0001111110100100";
                when "10100111" => z <= "0001111011110001";
                when "10101000" => z <= "0001111001000000";
                when "10101001" => z <= "0001110110010001";
                when "10101010" => z <= "0001110011100100";
                when "10101011" => z <= "0001110000111001";
                when "10101100" => z <= "0001101110010000";
                when "10101101" => z <= "0001101011101001";
                when "10101110" => z <= "0001101001000100";
                when "10101111" => z <= "0001100110100001";
                when "10110000" => z <= "0001100100000000";
                when "10110001" => z <= "0001100001100001";
                when "10110010" => z <= "0001011111000100";
                when "10110011" => z <= "0001011100101001";
                when "10110100" => z <= "0001011010010000";
                when "10110101" => z <= "0001010111111001";
                when "10110110" => z <= "0001010101100100";
                when "10110111" => z <= "0001010011010001";
                when "10111000" => z <= "0001010001000000";
                when "10111001" => z <= "0001001110110001";
                when "10111010" => z <= "0001001100100100";
                when "10111011" => z <= "0001001010011001";
                when "10111100" => z <= "0001001000010000";
                when "10111101" => z <= "0001000110001001";
                when "10111110" => z <= "0001000100000100";
                when "10111111" => z <= "0001000010000001";
                when "11000000" => z <= "0001000000000000";
                when "11000001" => z <= "0000111110000001";
                when "11000010" => z <= "0000111100000100";
                when "11000011" => z <= "0000111010001001";
                when "11000100" => z <= "0000111000010000";
                when "11000101" => z <= "0000110110011001";
                when "11000110" => z <= "0000110100100100";
                when "11000111" => z <= "0000110010110001";
                when "11001000" => z <= "0000110001000000";
                when "11001001" => z <= "0000101111010001";
                when "11001010" => z <= "0000101101100100";
                when "11001011" => z <= "0000101011111001";
                when "11001100" => z <= "0000101010010000";
                when "11001101" => z <= "0000101000101001";
                when "11001110" => z <= "0000100111000100";
                when "11001111" => z <= "0000100101100001";
                when "11010000" => z <= "0000100100000000";
                when "11010001" => z <= "0000100010100001";
                when "11010010" => z <= "0000100001000100";
                when "11010011" => z <= "0000011111101001";
                when "11010100" => z <= "0000011110010000";
                when "11010101" => z <= "0000011100111001";
                when "11010110" => z <= "0000011011100100";
                when "11010111" => z <= "0000011010010001";
                when "11011000" => z <= "0000011001000000";
                when "11011001" => z <= "0000010111110001";
                when "11011010" => z <= "0000010110100100";
                when "11011011" => z <= "0000010101011001";
                when "11011100" => z <= "0000010100010000";
                when "11011101" => z <= "0000010011001001";
                when "11011110" => z <= "0000010010000100";
                when "11011111" => z <= "0000010001000001";
                when "11100000" => z <= "0000010000000000";
                when "11100001" => z <= "0000001111000001";
                when "11100010" => z <= "0000001110000100";
                when "11100011" => z <= "0000001101001001";
                when "11100100" => z <= "0000001100010000";
                when "11100101" => z <= "0000001011011001";
                when "11100110" => z <= "0000001010100100";
                when "11100111" => z <= "0000001001110001";
                when "11101000" => z <= "0000001001000000";
                when "11101001" => z <= "0000001000010001";
                when "11101010" => z <= "0000000111100100";
                when "11101011" => z <= "0000000110111001";
                when "11101100" => z <= "0000000110010000";
                when "11101101" => z <= "0000000101101001";
                when "11101110" => z <= "0000000101000100";
                when "11101111" => z <= "0000000100100001";
                when "11110000" => z <= "0000000100000000";
                when "11110001" => z <= "0000000011100001";
                when "11110010" => z <= "0000000011000100";
                when "11110011" => z <= "0000000010101001";
                when "11110100" => z <= "0000000010010000";
                when "11110101" => z <= "0000000001111001";
                when "11110110" => z <= "0000000001100100";
                when "11110111" => z <= "0000000001010001";
                when "11111000" => z <= "0000000001000000";
                when "11111001" => z <= "0000000000110001";
                when "11111010" => z <= "0000000000100100";
                when "11111011" => z <= "0000000000011001";
                when "11111100" => z <= "0000000000010000";
                when "11111101" => z <= "0000000000001001";
                when "11111110" => z <= "0000000000000100";
                when "11111111" => z <= "0000000000000001";
                when others => z <= "0000000000000000";
            end case;
        end if;
    end process;
end rtl;
